

out clk;
